----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12.11.2024 09:24:03
-- Design Name: 
-- Module Name: SignalLatch - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SignalLatch is
 Port (
    clk_12M : in std_logic;
    drdy_in : in std_logic;
    drdy_latch : out std_logic
  );
end SignalLatch;

architecture Behavioral of SignalLatch is
    signal temp : std_logic := '0';
begin

    process (clk_12M, drdy_in)        
    begin
    
    if (rising_edge(drdy_in)) then
        drdy_latch <= '1';
        if(clk_12M = '1') then
            temp <= '1';        
        end if;
    end if;
          if (falling_edge(clk_12M)) then
        if(temp = '1') then
            temp <= '0';
        else
            drdy_latch <= '0';
        end if;
    end if;
   
    end process;
   


end Behavioral;
